`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.03.2023 12:59:47
// Design Name: 
// Module Name: find_the_white
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module find_the_white(
    input clock,
    input mouse_left_click,
    input [6:0] x, y,
    output reg [15:0] oled_data = 0
    );
    reg[95:0] r2 = 96'b011111101111110111111011001101100000110001111110110011011111100000111101100000011011111101111110;
    reg[95:0] r3 = 96'b011111101111110111111011001101100000110001111110110011011111100001111101100000011011111101111110;
    reg[95:0] r4 = 96'b000001100011000001100011001101100000110000000110110011000110000011101101100001111000110000000110;
    reg[95:0] r5 = 96'b000001100011000001100011001101100000110000000110110011000110000011001101100001111000110000000110;
    reg[95:0] r6 = 96'b011111100011000001100011111101101110110001111110111111000110000011001101100110011000110000011110;
    reg[95:0] r7 = 96'b011111100011000001100011111101101110110001111110111111000110000011001101100110011000110000011110;
    reg[95:0] r8 = 96'b000001100011000001100011001100111111100000000110110011000110000011001101111000011000110000000110;
    reg[95:0] r9 = 96'b000001100011000001100011001100111111100000000110110011000110000011101101111000011000110000000110;
    reg[95:0] r10 = 96'b011111100011000111111011001100011011000001111110110011000110000001111101100000011011111100000110;
    reg[95:0] r11 = 96'b011111100011000111111011001100011011000001111110110011000110000000111101100000011011111100000110;
    
    reg[95:0] r15 = 96'b000000000000000111100000000011110000011111111111111111111111000001111100000000000000000011111000;
    reg[95:0] r16 = 96'b000000000000000111100000000011110000011111111111111111111111000001111100000000000000000011111000;
    reg[95:0] r17 = 96'b000000000000000111100000000111110000011111111111111111111111000001111100000000000000000011111000;
    reg[95:0] r18 = 96'b000000000000000111100000000111110000011111111111111111111111000001111100000000000000000011111000;
    reg[95:0] r19 = 96'b000000000000000111100000001111110000000000000011111000000000000000111110000000000000000111110000;
    reg[95:0] r20 = 96'b000000000000000111100000001111110000000000000011111000000000000000111110000000000000000111110000;
    reg[95:0] r21 = 96'b000000000000000111100000011111110000000000000011111000000000000000011110000000000000000111100000;
    reg[95:0] r22 = 96'b000000000000000111100000011111110000000000000011111000000000000000011110000000000000000111100000;
    reg[95:0] r23 = 96'b000000000000000111100000111111110000000000000011111000000000000000011111000000000000001111100000;
    reg[95:0] r24 = 96'b000000000000000111100000111111110000000000000011111000000000000000011111000000000000001111100000;
    reg[95:0] r25 = 96'b000000000000000111100001111111110000000000000011111000000000000000001111000000000000001111000000;
    reg[95:0] r26 = 96'b000000000000000111100001111111110000000000000011111000000000000000001111000000000000001111000000;
    reg[95:0] r27 = 96'b000000000000000111100011111011110000000000000011111000000000000000001111100000000000011111000000;
    reg[95:0] r28 = 96'b000000000000000111100011111011110000000000000011111000000000000000001111100001111000011111000000;
    reg[95:0] r29 = 96'b000000000000000111100111110011110000000000000011111000000000000000000111100001111000011110000000;
    reg[95:0] r30 = 96'b000000000000000111100111110011110000000000000011111000000000000000000111100001111000011110000000;
    reg[95:0] r31 = 96'b000000000000000111101111100011110000000000000011111000000000000000000111110001111000111110000000;
    reg[95:0] r32 = 96'b000000000000000111101111100011110000000000000011111000000000000000000111110011111100111110000000;
    reg[95:0] r33 = 96'b000000000000000111111111000011110000000000000011111000000000000000000011111111111111111100000000;
    reg[95:0] r34 = 96'b000000000000000111111111000011110000000000000011111000000000000000000011111111111111111100000000;
    reg[95:0] r35 = 96'b000000000000000111111110000011110000000000000011111000000000000000000011111111111111111100000000;
    reg[95:0] r36 = 96'b000000000000000111111110000011110000000000000011111000000000000000000011111111111111111100000000;
    reg[95:0] r37 = 96'b000000000000000111111100000011110000000000000011111000000000000000000001111111111111111000000000;
    reg[95:0] r38 = 96'b000000000000000111111100000011110000000000000011111000000000000000000001111111111111111000000000;
    reg[95:0] r39 = 96'b000000000000000111111000000011110000000000000011111000000000000000000001111111111111111000000000;
    reg[95:0] r40 = 96'b000000000000000111111000000011110000011111111111111111111111000000000001111111001111111000000000;
    reg[95:0] r41 = 96'b000000000000000111110000000011110000011111111111111111111111000000000000111111001111110000000000;
    reg[95:0] r42 = 96'b000000000000000111110000000011110000011111111111111111111111000000000000111111001111110000000000;
    reg[95:0] r43 = 96'b000000000000000111100000000011110000011111111111111111111111000000000000111111001111110000000000;
    
    reg [15:0] color_hex = 0;
    
    always @(posedge clock)
    begin
        color_hex <= mouse_left_click ? color_hex + 1 : color_hex ;
        if ((y == 2 && r2[x]==1) || (y == 3 && r3[x]==1) || (y == 4 && r4[x]==1) || (y == 5 && r5[x]==1)
         || (y == 6 && r6[x]==1) || (y == 7 && r7[x]==1) || (y == 8 && r8[x]==1) || (y == 9 && r9[x]==1)
         || (y == 10 && r10[x]==1) || (y == 11 && r11[x]==1))
        begin
            oled_data <= 16'hffff;
        end
        else
        begin
            if (color_hex <= 16'hffff && color_hex >= 16'hfdef)
            begin
                if ((y == 15 && r15[x]==1) || (y == 16 && r16[x]==1) || (y == 17 && r17[x]==1) 
                || (y == 18 && r18[x]==1) || (y == 19 && r19[x]==1) || (y == 20 && r20[x]==1) 
                || (y == 21 && r21[x]==1) || (y == 22 && r22[x]==1) || (y == 23 && r23[x]==1) 
                || (y == 24 && r24[x]==1) || (y == 25 && r25[x]==1) || (y == 26 && r26[x]==1) 
                || (y == 27 && r27[x]==1) || (y == 28 && r28[x]==1) || (y == 29 && r29[x]==1) 
                || (y == 30 && r30[x]==1) || (y == 31 && r31[x]==1) || (y == 32 && r32[x]==1) 
                || (y == 33 && r33[x]==1) || (y == 34 && r34[x]==1) || (y == 35 && r35[x]==1) 
                || (y == 36 && r36[x]==1) || (y == 37 && r37[x]==1) || (y == 38 && r38[x]==1) 
                || (y == 39 && r39[x]==1) || (y == 40 && r40[x]==1) || (y == 41 && r41[x]==1) 
                || (y == 42 && r42[x]==1) || (y == 43 && r43[x]==1))
                begin
                    oled_data <= 0;
                end
                else 
                begin
                    oled_data <= 16'hffff;
                end
            end
            else
            begin
                oled_data <= color_hex;              
            end
        end
    end
endmodule
